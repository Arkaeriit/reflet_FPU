../floating_points_operations/reflet_float_functions.vh