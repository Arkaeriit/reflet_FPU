/*----------------------------------------\
|This file contains constants used by some|
|floating point opperations. The value of |
|the multiplier time should be changed    |
|depending on the integer multiplier used.|
\----------------------------------------*/

`ifndef reflet_float_opperations
`define reflet_float_opperations

`define multiplication_time 2

`endif

