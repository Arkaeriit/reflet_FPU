../float_processing/reflet_fpu.vh